library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

package CONSTANTS is
   constant N: integer := 32;
end package;

	


